module help

pub fn show_help() {
    println('lana - Vlang C++ Build System')
    println('Usage: lana [command] [options]')
    println('')
    println('Commands:')
    println('  build           Build the project')
    println('  clean           Clean build files')
    println('  run             Build and run the project')
    println('  init <name>     Initialize new project')
    println('')
    println('Options:')
    println('  -d, --debug     Enable debug mode')
    println('  -O, --optimize  Enable optimization')
    println('  -v, --verbose   Verbose output')
    println('  -o, --output    Set output name')
    println('  -I <dir>        Add include directory')
    println('  -l <lib>        Add library')
    println('  --config <file> Use config file')
    println('')
    println('Examples:')
    println('  lana build -d -I include/mylib')
    println('  lana run')
    println('  lana init myproject')
    println('')
    println('Project Structure:')
    println('  src/      - Source files (.cpp, .cc, .cxx)')
    println('  include/  - Header files (.h, .hpp)')
    println('  build/    - Object files and intermediates')
    println('  bin/      - Executable output')
    println('  config.ini - Build configuration')
}