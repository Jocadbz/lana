module help

pub fn show_help() {
    println('lana - Vlang C++ Build System')
    println('Usage: lana [command] [options]')
    println('')
    println('Commands:')
    println('  build           Build the project (shared libs + tools)')
    println('  clean           Clean build files')
    println('  run             Build and run the main tool')
    println('  init <name>     Initialize new project')
    println('')
    println('Options:')
    println('  -d, --debug     Enable debug mode')
    println('  -O, --optimize  Enable optimization')
    println('  -v, --verbose   Verbose output')
    println('  -p, --parallel  Enable parallel compilation')
    println('  -o, --output    Set output name')
    println('  -I <dir>        Add include directory')
    println('  -l <lib>        Add library')
    println('  --config <file> Use config file')
    println('  --shared-lib <name> <source>  Add shared library')
    println('  --tool <name> <source>        Add tool/executable')
    println('')
    println('Configuration File (config.ini):')
    println('  [global]')
    println('  project_name = myproject')
    println('  src_dir = src')
    println('  debug = true')
    println('  ')
    println('  [shared_libs]')
    println('  name = net')
    println('  sources = src/lib/net/connection.cpp')
    println('  libraries = cli')
    println('  ')
    println('  [tools]')
    println('  name = dumpnbt')
    println('  sources = src/tools/dumpnbt.cpp')
    println('  libraries = nbt,cli')
    println('')
    println('Examples:')
    println('  lana build -d -v -p')
    println('  lana run')
    println('  lana build --shared-lib cli src/lib/cli.cpp --tool dumpnbt src/tools/dumpnbt.cpp')
    println('  lana init myproject')
    println('')
    println('Project Structure:')
    println('  src/           - Source files (.cpp, .cc, .cxx)')
    println('    lib/         - Shared library sources')
    println('    tools/       - Tool/executable sources')
    println('  include/       - Header files (.h, .hpp)')
    println('  build/         - Object files and intermediates')
    println('  bin/           - Output')
    println('    lib/         - Shared libraries (.so/.dll)')
    println('    tools/       - Executables')
    println('  config.ini     - Build configuration')
}