module help

import docstore

pub fn show_help() {
    print(docstore.help_text())
}